--Simple Counter
