library verilog;
use verilog.vl_types.all;
entity Flancter_vlg_vec_tst is
end Flancter_vlg_vec_tst;
