library verilog;
use verilog.vl_types.all;
entity testing_top_vlg_vec_tst is
end testing_top_vlg_vec_tst;
